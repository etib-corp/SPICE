boolean: ["true", "false"]
variable{suffix: ";"}: ["let", "const", "var"]
operators{suffix: ";"}: [plus: expression -> "+" -> expression, minus: expression -> "-" -> expression, multiply: expression -> "*" -> expression, divide: expression -> "/" -> expression, modulo: expression -> "%" -> expression, equal: expression -> ["==", "==="] -> expression, assignation: name -> "=" -> expression]
condition{prefix: "(", suffix: ")"}: expression
parameters{prefix: "(", suffix: ")"}: name -> ","
codeBlock{prefix: "{", suffix: "}"}: many(expression)
if: ["if"] -> condition -> codeBlock
function: ["function"] -> name -> parameters -> codeBlock