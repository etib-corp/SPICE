boolean{prefix: "(", suffix: ")"}: ["#t", "#f"]
variable{prefix: "(", suffix: ")"}: ["define"]
operators{prefix: "(", suffix: ")"}: [plus: "+" -> expression -> expression, minus: "-" -> expression -> expression, multiply: "*" -> expression -> expression, divide: "/" -> expression -> expression, modulo: "%" -> expression -> expression, equal: "eq?" -> expression -> expression, assignation: name -> "=" -> expression]
condition{prefix: "(", suffix: ")"}: expression
parameters{prefix: "(", suffix: ")"}: name -> " "
codeBlock{prefix: "(", suffix: ")"}: ["\n"]
if{prefix: "(", suffix: ")"}: ["if"] -> [""]
function{prefix: "(", suffix: ")"}: ["define"] -> name -> parameters -> codeBlock
