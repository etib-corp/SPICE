boolean{prefix:"(", suffix:")"}: ["true", "false"]
variable{prefix:"", suffix: ""}: ["let", "const", "var"]
operators: [plus: expression -> "+" -> expression , minus: expression -> "-" -> expression , multiply: expression -> "*" -> expression , divide: expression -> "/" -> expression , modulo: expression -> "%" -> expression , equal: expression -> "===" -> expression , assignation: expression -> "=" -> expression, less: expression -> "<" -> expression, greater: expression -> ">" -> expression]
condition{prefix: "(", suffix: ")"}: expression
parameters{prefix: "(", suffix: ")"}: name -> ","
codeBlock{prefix: "{", suffix: "}"}: [";"]
if: ["if"] -> ["else"]
function: ["function"] -> name -> parameters -> codeBlock
